
interface intf(input bit clk);
    // ------------------- port declaration-------------------------------------
    logic [7:0]in1;
    logic [7:0]in2;
    logic [15:0]out;

endinterface

